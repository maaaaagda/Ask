CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 110 17 150 10
176 80 1364 520
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 2 0.283892 0.500000
176 529 1364 707
42991634 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 378 343 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89562e-315 0
0
13 Logic Switch~
5 43 175 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-4 -30 10 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89562e-315 0
0
9 Inverter~
13 105 277 0 2 22
0 2 12
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U8A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3124 0 0
2
42473.7 0
0
5 4001~
219 530 253 0 3 22
0 7 6 13
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
3421 0 0
2
42473.7 0
0
5 4001~
219 529 205 0 3 22
0 5 8 14
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
8157 0 0
2
42473.7 0
0
5 4011~
219 223 269 0 3 22
0 5 12 11
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
5572 0 0
2
42473.7 0
0
5 4011~
219 305 211 0 3 22
0 10 11 9
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
8901 0 0
2
42473.7 0
0
5 4011~
219 234 165 0 3 22
0 6 2 10
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
7361 0 0
2
42473.7 0
0
5 SCOPE
12 379 273 0 1 11
0 3
0
0 0 57584 0
3 TP4
-11 -4 10 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4747 0 0
2
42473.6 0
0
5 SCOPE
12 125 165 0 1 11
0 2
0
0 0 57584 0
3 TP3
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
972 0 0
2
42473.6 0
0
5 SCOPE
12 591 182 0 1 11
0 13
0
0 0 57584 0
3 TP2
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3472 0 0
2
42473.6 0
0
5 SCOPE
12 570 182 0 1 11
0 14
0
0 0 57584 0
3 TP1
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9998 0 0
2
42473.6 0
0
2 +V
167 308 283 0 1 3
0 3
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
5.89562e-315 0
0
14 Logic Display~
6 593 157 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.89562e-315 0
0
14 Logic Display~
6 570 158 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.89562e-315 0
0
6 74LS74
17 454 233 0 12 25
0 4 9 3 3 4 5 3 3 5
6 7 8
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.89562e-315 0
0
27
1 0 2 0 0 4096 0 10 0 0 19 2
125 177
125 175
1 0 3 0 0 0 0 9 0 0 3 2
379 285
379 285
8 0 3 0 0 8192 0 16 0 0 4 3
416 269
416 285
353 285
0 1 3 0 0 8320 0 0 13 25 0 5
416 219
353 219
353 296
308 296
308 292
5 0 4 0 0 4096 0 16 0 0 6 2
422 242
403 242
1 1 4 0 0 8320 0 16 1 0 0 4
422 197
403 197
403 343
390 343
0 1 5 0 0 4096 0 0 5 9 0 4
486 182
511 182
511 196
516 196
0 1 6 0 0 8320 0 0 8 11 0 5
492 224
492 127
187 127
187 156
210 156
9 0 5 0 0 8192 0 16 0 0 10 4
486 206
486 151
341 151
341 251
1 6 5 0 0 12416 0 6 16 0 0 4
199 260
178 260
178 251
422 251
10 2 6 0 0 0 0 16 4 0 0 4
492 215
492 233
517 233
517 262
11 1 7 0 0 12416 0 16 4 0 0 4
486 251
492 251
492 244
517 244
12 2 8 0 0 8320 0 16 5 0 0 4
492 260
499 260
499 214
516 214
3 2 9 0 0 12416 0 7 16 0 0 4
332 211
372 211
372 206
422 206
3 1 10 0 0 4224 0 8 7 0 0 3
261 165
261 202
281 202
3 2 11 0 0 8320 0 6 7 0 0 4
250 269
265 269
265 220
281 220
2 2 12 0 0 8320 0 3 6 0 0 3
126 277
126 278
199 278
0 1 2 0 0 4096 0 0 3 19 0 3
60 175
60 277
90 277
1 2 2 0 0 4224 0 2 8 0 0 4
55 175
201 175
201 174
210 174
3 0 13 0 0 4096 0 4 0 0 26 2
569 253
569 254
3 0 14 0 0 4096 0 5 0 0 27 2
568 205
570 205
1 0 13 0 0 0 0 11 0 0 26 2
591 194
592 194
1 0 14 0 0 0 0 12 0 0 27 2
570 194
570 194
7 8 3 0 0 0 0 16 16 0 0 2
416 260
416 269
3 4 3 0 0 0 0 16 16 0 0 2
416 215
416 224
0 1 13 0 0 8320 0 0 14 0 0 4
566 254
592 254
592 175
593 175
1 0 14 0 0 4224 0 15 0 0 0 3
570 176
570 206
565 206
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
