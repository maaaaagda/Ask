CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 311 319 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
42474.9 0
0
13 Logic Switch~
5 286 231 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
42474.9 1
0
5 4001~
219 605 250 0 3 22
0 6 9 5
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
3124 0 0
2
42474.9 0
0
5 4001~
219 584 338 0 3 22
0 6 8 7
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
3421 0 0
2
42474.9 0
0
6 74LS76
104 470 263 0 14 29
0 4 4 2 3 3 10 11 12 13
14 9 8 15 16
0
0 0 4848 0
6 74LS76
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=13;
130 %D [%5bi %13bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 16 1 2 3 9 12 6 7
8 15 14 11 10 4 16 1 2 3
9 12 6 7 8 15 14 11 10 0
65 0 0 512 0 0 0 0
1 U
8157 0 0
2
42474.9 0
0
2 +V
167 288 341 0 1 3
0 3
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
5.89657e-315 0
0
14 Logic Display~
6 656 334 0 1 2
10 7
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
42474.9 2
0
14 Logic Display~
6 692 247 0 1 2
10 5
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
42474.9 3
0
9 Inverter~
13 546 241 0 2 22
0 4 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4747 0 0
2
42474.9 7
0
14
3 1 2 0 0 4224 0 5 1 0 0 4
432 245
329 245
329 319
323 319
0 0 3 0 0 4096 0 0 0 4 3 2
392 263
342 263
4 1 3 0 0 8320 0 5 6 0 0 4
432 254
342 254
342 350
288 350
5 0 3 0 0 0 0 5 0 0 0 2
432 263
388 263
0 5 3 0 0 0 0 0 5 0 0 2
438 263
432 263
1 0 4 0 0 4096 0 2 0 0 7 4
298 231
343 231
343 227
358 227
0 2 4 0 0 8192 0 0 5 8 0 3
358 227
358 236
438 236
1 1 4 0 0 8320 0 9 5 0 0 5
531 241
531 186
358 186
358 227
438 227
3 1 5 0 0 8320 0 3 8 0 0 3
644 250
644 251
676 251
2 1 6 0 0 4096 0 9 3 0 0 2
567 241
592 241
3 1 7 0 0 4224 0 4 7 0 0 2
623 338
640 338
12 2 8 0 0 12416 0 5 4 0 0 5
508 236
508 276
528 276
528 347
571 347
11 2 9 0 0 12416 0 5 3 0 0 4
502 227
519 227
519 259
592 259
2 1 6 0 0 4224 0 9 4 0 0 5
567 241
567 303
553 303
553 329
571 329
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
