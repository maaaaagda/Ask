CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
410 0 1 200 10
184 87 673 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
13 C:\CM\BOM.DAT
0 7
5 4 0.235825 0.500000
352 183 465 280
177209362 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 171 284 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
1 d
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
41729.3 0
0
13 Logic Switch~
5 170 232 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -17 8 -9
1 c
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
41729.3 1
0
13 Logic Switch~
5 171 177 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
1 b
-4 -27 3 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
41729.3 2
0
13 Logic Switch~
5 169 122 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21088 0
2 5V
-6 -16 8 -8
1 a
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
41729.3 3
0
2 +V
167 489 255 0 1 3
0 2
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.8956e-315 0
0
14 Logic Display~
6 577 150 0 1 2
10 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
41729.3 4
0
6 74LS74
17 505 195 0 12 25
0 5 4 2 2 14 15 16 17 3
4 18 19
0
0 0 4832 0
6 74LS74
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 512 1 0 0 0
1 U
8901 0 0
2
41729.3 5
0
5 4023~
219 309 179 0 4 22
0 8 7 6 9
0
0 0 608 0
4 4023
-14 -28 14 -20
6 NAND3A
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 1 2 0
1 U
7361 0 0
2
5.8956e-315 5.26354e-315
0
5 4023~
219 395 194 0 4 22
0 13 9 12 5
0
0 0 608 0
4 4023
-14 -28 14 -20
6 NAND3C
-21 -25 21 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 3 4 0
1 U
4747 0 0
2
5.8956e-315 5.30499e-315
0
10 2-In NAND~
219 315 131 0 3 22
0 11 6 13
0
0 0 608 0
4 4011
-7 -24 21 -16
5 NAND2
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 5 0
1 U
972 0 0
2
5.8956e-315 5.32571e-315
0
5 4023~
219 291 235 0 4 22
0 8 7 10 12
0
0 0 608 0
4 4023
-14 -28 14 -20
6 NAND3B
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 2 0
65 0 0 0 3 2 4 0
1 U
3472 0 0
2
5.8956e-315 5.34643e-315
0
9 Inverter~
13 221 122 0 2 22
0 10 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 1 0
1 U
9998 0 0
2
41729.3 6
0
14 Logic Display~
6 443 241 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
41729.3 7
0
20
8 0 0 0 0 0 0 7 0 0 3 2
467 231
467 231
7 0 0 0 0 0 0 7 0 0 3 2
467 222
467 222
4 1 2 0 0 4224 0 7 5 0 0 3
467 186
467 264
489 264
3 4 2 0 0 0 0 7 7 0 0 2
467 177
467 186
9 1 3 0 0 8320 0 7 6 0 0 4
537 168
549 168
549 154
561 154
2 10 4 0 0 12416 0 7 7 0 0 6
473 168
463 168
463 125
551 125
551 177
543 177
1 0 5 0 0 8320 0 7 0 0 8 4
473 159
448 159
448 195
443 195
1 4 5 0 0 0 0 13 9 0 0 3
443 227
443 194
422 194
0 3 6 0 0 4096 0 0 8 18 0 2
226 188
285 188
0 2 7 0 0 4096 0 0 8 14 0 3
240 232
240 179
285 179
1 1 8 0 0 8320 0 3 8 0 0 3
183 177
183 170
285 170
4 2 9 0 0 8320 0 8 9 0 0 3
336 179
336 194
371 194
0 3 10 0 0 4224 0 0 11 17 0 3
194 122
194 244
267 244
1 2 7 0 0 4224 0 2 11 0 0 4
182 232
259 232
259 235
267 235
1 1 8 0 0 0 0 3 11 0 0 5
183 177
183 204
259 204
259 226
267 226
2 1 11 0 0 4224 0 12 10 0 0 2
242 122
291 122
1 1 10 0 0 0 0 4 12 0 0 2
181 122
206 122
1 2 6 0 0 8320 0 1 10 0 0 4
183 284
226 284
226 140
291 140
4 3 12 0 0 4224 0 11 9 0 0 4
318 235
357 235
357 203
371 203
1 3 13 0 0 8320 0 9 10 0 0 4
371 185
357 185
357 131
342 131
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
