CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 79 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 357 256 0 1 11
0 8
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89606e-315 0
0
13 Logic Switch~
5 360 178 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89606e-315 5.26354e-315
0
13 Logic Switch~
5 357 219 0 1 11
0 7
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89606e-315 5.30499e-315
0
14 Logic Display~
6 547 329 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L4
-7 25 7 33
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.89606e-315 5.32571e-315
0
14 Logic Display~
6 624 329 0 1 2
10 3
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
-9 23 5 31
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89606e-315 5.34643e-315
0
14 Logic Display~
6 600 329 0 1 2
10 4
0
0 0 53872 692
6 100MEG
3 -16 45 -8
2 L2
-7 24 7 32
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89606e-315 5.3568e-315
0
14 Logic Display~
6 573 329 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
-7 25 7 33
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89606e-315 5.36716e-315
0
7 Ground~
168 538 229 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
5.89606e-315 5.37752e-315
0
7 74LS194
49 470 234 0 14 29
0 9 7 8 10 6 7 7 2 2
2 3 4 5 6
0
0 0 4832 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.89606e-315 5.38788e-315
0
13
11 1 3 0 0 4224 0 9 5 0 0 3
502 243
624 243
624 315
1 12 4 0 0 8320 0 6 9 0 0 3
600 315
600 252
502 252
13 1 5 0 0 4224 0 9 7 0 0 3
502 261
573 261
573 315
0 1 6 0 0 4096 0 0 4 9 0 3
502 289
547 289
547 315
0 1 7 0 0 4096 0 0 3 6 0 2
404 219
369 219
0 7 7 0 0 8320 0 0 9 13 0 5
404 219
404 162
513 162
513 198
502 198
1 3 8 0 0 8320 0 1 9 0 0 5
369 256
369 237
439 237
439 225
438 225
1 1 9 0 0 8320 0 2 9 0 0 4
372 178
372 187
438 187
438 198
5 14 6 0 0 12416 0 9 9 0 0 5
438 252
432 252
432 289
502 289
502 270
0 1 2 0 0 4224 0 0 8 11 0 3
515 219
538 219
538 223
0 10 2 0 0 0 0 0 9 12 0 3
515 219
515 225
502 225
8 9 2 0 0 0 0 9 9 0 0 6
502 207
515 207
515 219
515 219
515 216
502 216
2 6 7 0 0 0 0 9 9 0 0 4
438 216
404 216
404 270
432 270
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
