CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 0 30 200 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 264 212 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
40983.5 0
0
13 Logic Switch~
5 297 131 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
40983.5 1
0
14 Logic Display~
6 617 84 0 1 2
12 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3124 0 0
2
40983.5 0
0
14 Logic Display~
6 596 84 0 1 2
21 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
40983.5 0
0
5 4001~
219 635 214 0 3 22
0 9 10 8
0
0 0 624 0
4 4001
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 4 0
1 U
8157 0 0
2
40983.5 2
0
5 4011~
219 441 192 0 3 22
0 14 7 4
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
40983.5 3
0
5 4011~
219 447 239 0 3 22
0 7 6 5
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 2 0
1 U
8901 0 0
2
40983.5 4
0
5 4011~
219 312 248 0 3 22
0 11 3 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 2 0
1 U
7361 0 0
2
40983.5 5
0
5 4011~
219 375 221 0 3 22
0 11 2 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
40983.5 6
0
5 4011~
219 370 183 0 3 22
0 9 11 14
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
40983.5 7
0
2 +V
167 451 99 0 1 3
0 13
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
40983.5 8
0
14 Logic Display~
6 659 145 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
40983.5 9
0
6 74LS74
17 531 187 0 12 25
0 12 4 13 13 12 5 13 13 3
9 2 10
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
40983.5 10
0
24
1 0 2 0 0 4096 0 3 0 0 8 4
617 102
617 190
569 190
569 205
1 0 3 0 0 4096 0 4 0 0 21 2
596 102
596 146
2 3 4 0 0 8320 0 13 6 0 0 3
499 160
468 160
468 192
6 3 5 0 0 8320 0 13 7 0 0 4
499 205
477 205
477 239
474 239
2 3 6 0 0 4224 0 7 8 0 0 2
423 248
339 248
0 1 7 0 0 4096 0 0 7 7 0 3
417 221
417 230
423 230
3 2 7 0 0 8320 0 9 6 0 0 3
402 221
417 221
417 201
2 11 2 0 0 8320 0 9 13 0 0 5
351 230
351 265
583 265
583 205
563 205
3 1 8 0 0 4224 0 5 12 0 0 3
674 214
674 163
659 163
1 10 9 0 0 12288 0 5 13 0 0 4
622 205
613 205
613 169
569 169
12 2 10 0 0 4224 0 13 5 0 0 4
569 214
609 214
609 223
622 223
1 0 11 0 0 4096 0 1 0 0 13 4
276 212
287 212
287 212
283 212
1 0 11 0 0 8192 0 8 0 0 23 3
288 239
283 239
283 212
5 0 12 0 0 8192 0 13 0 0 19 3
499 196
481 196
481 151
8 1 13 0 0 4224 0 13 11 0 0 3
493 223
493 108
451 108
7 8 13 0 0 0 0 13 13 0 0 2
493 214
493 223
4 7 13 0 0 0 0 13 13 0 0 2
493 178
493 214
3 4 13 0 0 0 0 13 13 0 0 2
493 169
493 178
1 1 12 0 0 12416 0 13 2 0 0 4
499 151
481 151
481 131
309 131
0 1 12 0 0 0 0 0 13 0 0 3
505 152
505 151
499 151
9 2 3 0 0 16512 0 13 8 0 0 7
563 160
563 146
598 146
598 275
276 275
276 257
288 257
10 1 9 0 0 12416 0 13 10 0 0 5
569 169
578 169
578 118
346 118
346 174
2 1 11 0 0 12416 0 10 9 0 0 4
346 192
283 192
283 212
351 212
3 1 14 0 0 4224 0 10 6 0 0 2
397 183
417 183
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
