CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 10 30 150 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 353 282 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
40988.4 0
0
13 Logic Switch~
5 353 242 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-4 -29 10 -21
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
40988.4 0
0
2 +V
167 308 283 0 1 3
0 2
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
40988.4 0
0
5 4081~
219 545 254 0 3 22
0 5 7 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3421 0 0
2
40988.4 0
0
5 4081~
219 544 206 0 3 22
0 6 7 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
8157 0 0
2
40988.4 0
0
14 Logic Display~
6 593 157 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5572 0 0
2
40988.4 0
0
14 Logic Display~
6 570 158 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
40988.4 0
0
6 74LS74
17 454 233 0 12 25
0 10 11 2 2 10 9 2 2 5
6 7 8
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 0 0 0 0 0
1 U
7361 0 0
2
40988.4 0
0
5 4071~
219 354 186 0 3 22
0 13 12 11
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
4747 0 0
2
40988.4 0
0
5 4081~
219 310 205 0 3 22
0 5 8 12
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1B
-13 -26 8 -18
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
972 0 0
2
40988.4 0
0
5 4081~
219 309 158 0 3 22
0 6 7 13
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
40988.4 0
0
20
8 1 2 0 0 8320 0 8 3 0 0 3
416 269
416 292
308 292
7 8 2 0 0 0 0 8 8 0 0 2
416 260
416 269
4 7 2 0 0 0 0 8 8 0 0 2
416 224
416 260
3 4 2 0 0 0 0 8 8 0 0 2
416 215
416 224
3 1 3 0 0 8336 0 4 6 0 0 4
566 254
592 254
592 175
593 175
1 3 4 0 0 4224 0 7 5 0 0 3
570 176
570 206
565 206
0 1 5 0 0 8320 0 0 10 8 0 5
502 245
502 316
274 316
274 196
286 196
9 1 5 0 0 0 0 8 4 0 0 4
486 206
494 206
494 245
521 245
0 1 6 0 0 8320 0 0 11 10 0 5
499 198
499 126
247 126
247 149
285 149
10 1 6 0 0 0 0 8 5 0 0 4
492 215
499 215
499 197
520 197
0 2 7 0 0 8320 0 0 11 12 0 5
512 215
512 112
238 112
238 167
285 167
0 2 7 0 0 0 0 0 5 13 0 3
512 251
512 215
520 215
11 2 7 0 0 0 0 8 4 0 0 4
486 251
512 251
512 263
521 263
12 2 8 0 0 8320 0 8 10 0 0 5
492 260
492 305
283 305
283 214
286 214
6 1 9 0 0 4224 0 8 2 0 0 3
422 251
365 251
365 242
1 0 10 0 0 8320 0 1 0 0 17 3
365 282
399 282
399 242
1 5 10 0 0 8320 0 8 8 0 0 4
422 197
399 197
399 242
422 242
2 3 11 0 0 4224 0 8 9 0 0 3
422 206
387 206
387 186
2 3 12 0 0 8320 0 9 10 0 0 4
341 195
336 195
336 205
331 205
3 1 13 0 0 8320 0 11 9 0 0 4
330 158
337 158
337 177
341 177
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
