CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 120 10
176 77 1278 749
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 173 457 270
42991634 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 311 319 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89657e-315 0
0
13 Logic Switch~
5 344 301 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89657e-315 0
0
2 +V
167 288 341 0 1 3
0 2
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
41736.1 0
0
10 2-In NAND~
219 547 338 0 3 22
0 11 8 4
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U6B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3421 0 0
2
41736.1 0
0
9 Inverter~
13 597 338 0 2 22
0 4 6
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8157 0 0
2
41736.1 0
0
10 2-In NAND~
219 543 241 0 3 22
0 12 8 5
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
5572 0 0
2
41736.1 0
0
14 Logic Display~
6 656 334 0 1 2
10 6
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89657e-315 0
0
14 Logic Display~
6 656 237 0 1 2
10 7
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.89657e-315 0
0
10 2-In NAND~
219 344 254 0 3 22
0 15 14 10
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
4747 0 0
2
5.89657e-315 0
0
10 2-In NAND~
219 295 272 0 3 22
0 11 13 14
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
972 0 0
2
5.89657e-315 0
0
10 2-In NAND~
219 283 221 0 3 22
0 12 8 15
0
0 0 624 0
6 74LS37
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3472 0 0
2
5.89657e-315 0
0
9 Inverter~
13 593 241 0 2 22
0 5 7
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9998 0 0
2
5.89657e-315 0
0
6 74LS74
17 432 282 0 12 25
0 9 10 2 2 9 3 2 2 11
12 8 13
0
0 0 4848 0
6 74LS74
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 0
65 0 0 0 1 0 0 0
1 U
3536 0 0
2
5.89657e-315 0
0
22
8 0 2 0 0 4096 0 13 0 0 2 2
394 318
386 318
1 3 2 0 0 8320 0 3 13 0 0 5
288 350
288 348
386 348
386 264
394 264
6 1 3 0 0 8320 0 13 2 0 0 3
400 300
400 301
356 301
3 1 4 0 0 4224 0 4 5 0 0 2
574 338
582 338
3 1 5 0 0 4224 0 6 12 0 0 2
570 241
578 241
2 1 6 0 0 4224 0 5 7 0 0 2
618 338
640 338
2 1 7 0 0 4224 0 12 8 0 0 2
614 241
640 241
11 0 8 0 0 4096 0 13 0 0 20 2
464 300
492 300
5 0 9 0 0 4096 0 13 0 0 10 2
400 291
371 291
1 1 9 0 0 8320 0 13 1 0 0 5
400 246
371 246
371 320
323 320
323 319
2 3 10 0 0 8320 0 13 9 0 0 3
400 255
400 254
371 254
2 0 8 0 0 0 0 6 0 0 20 2
519 250
492 250
7 0 2 0 0 0 0 13 0 0 2 2
394 309
386 309
0 4 2 0 0 0 0 0 13 2 0 4
386 272
383 272
383 273
394 273
0 1 11 0 0 4096 0 0 4 16 0 2
502 329
523 329
1 9 11 0 0 12416 0 10 13 0 0 6
271 263
227 263
227 370
502 370
502 255
464 255
1 0 12 0 0 4096 0 6 0 0 18 2
519 232
478 232
1 10 12 0 0 12416 0 11 13 0 0 6
259 212
257 212
257 181
478 181
478 264
470 264
2 12 13 0 0 12416 0 10 13 0 0 6
271 281
241 281
241 358
477 358
477 309
470 309
2 2 8 0 0 12416 0 11 4 0 0 6
259 230
242 230
242 168
492 168
492 347
523 347
2 3 14 0 0 4224 0 9 10 0 0 3
320 263
320 272
322 272
1 3 15 0 0 8320 0 9 11 0 0 3
320 245
310 245
310 221
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
