CircuitMaker Text
5.6
Probes: 1
v1[p]
Operating Point
0 294 341 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 210 30 200 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 450 266 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89559e-315 0
0
13 Logic Switch~
5 415 338 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89559e-315 5.26354e-315
0
10 3-In NAND~
219 575 366 0 4 22
0 8 7 6 5
0
0 0 624 0
5 74F10
-18 -28 17 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
3124 0 0
2
5.89559e-315 5.30499e-315
0
7 Ground~
168 453 301 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
5.89559e-315 5.32571e-315
0
14 Logic Display~
6 557 270 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.89559e-315 5.34643e-315
0
14 Logic Display~
6 578 270 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89559e-315 5.3568e-315
0
14 Logic Display~
6 599 270 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89559e-315 5.36716e-315
0
14 Logic Display~
6 621 269 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.89559e-315 5.37752e-315
0
7 74LS194
49 497 302 0 14 29
0 3 4 2 10 5 4 11 12 13
14 8 7 6 9
0
0 0 4848 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.89559e-315 5.38788e-315
0
12
1 1 3 0 0 4224 0 1 9 0 0 2
462 266
465 266
1 0 4 0 0 4096 0 2 0 0 3 2
427 338
435 338
2 6 4 0 0 8320 0 9 9 0 0 4
465 284
435 284
435 338
459 338
5 4 5 0 0 12416 0 9 3 0 0 6
465 320
456 320
456 388
606 388
606 366
602 366
3 0 6 0 0 8192 0 3 0 0 8 3
551 375
530 375
530 329
0 2 7 0 0 4096 0 0 3 10 0 3
538 320
538 366
551 366
0 1 8 0 0 4224 0 0 3 11 0 3
547 311
547 357
551 357
13 1 6 0 0 4224 0 9 7 0 0 3
529 329
599 329
599 288
1 3 2 0 0 8320 0 4 9 0 0 3
453 295
453 293
465 293
1 12 7 0 0 8320 0 6 9 0 0 3
578 288
578 320
529 320
11 1 8 0 0 0 0 9 5 0 0 3
529 311
557 311
557 288
14 1 9 0 0 4224 0 9 8 0 0 3
529 338
621 338
621 287
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
