CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 160 1 210 10
176 79 1364 558
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 1 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 2 0.235110 0.500000
176 567 1364 717
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 385 285 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 RES
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
5.89467e-315 0
0
5 SCOPE
12 708 187 0 1 11
0 3
0
0 0 57584 0
2 Q0
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6357 0 0
2
40240.6 0
0
5 SCOPE
12 671 188 0 1 11
0 4
0
0 0 57584 0
2 Q1
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
319 0 0
2
40240.6 0
0
5 SCOPE
12 636 188 0 1 11
0 5
0
0 0 57584 0
2 Q2
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3976 0 0
2
40240.6 0
0
5 SCOPE
12 600 188 0 1 11
0 6
0
0 0 57584 0
2 Q3
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7634 0 0
2
40240.6 0
0
5 SCOPE
12 293 191 0 1 11
0 7
0
0 0 57584 0
3 RES
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
523 0 0
2
40240.6 0
0
5 SCOPE
12 372 191 0 1 11
0 8
0
0 0 57584 0
3 CLK
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6748 0 0
2
40240.6 0
0
7 Pulser~
4 329 267 0 10 12
0 10 11 8 12 0 0 2 2 2
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6901 0 0
2
5.89467e-315 5.26354e-315
0
14 Logic Display~
6 575 230 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
5.89467e-315 5.38788e-315
0
14 Logic Display~
6 555 230 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
5.89467e-315 5.39306e-315
0
14 Logic Display~
6 534 230 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
5.89467e-315 5.39824e-315
0
14 Logic Display~
6 513 230 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
5.89467e-315 5.40342e-315
0
7 Ground~
168 500 376 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5551 0 0
2
5.89467e-315 5.4086e-315
0
2 +V
167 406 217 0 1 3
0 9
0
0 0 54256 0
2 5V
-8 -22 6 -14
3 VCC
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6986 0 0
2
5.89467e-315 5.41378e-315
0
7 74LS194
49 449 294 0 14 29
0 8 9 7 13 3 9 9 2 2
2 6 5 4 3
0
0 0 4848 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
8745 0 0
2
5.89467e-315 5.41896e-315
0
19
1 0 3 0 0 8336 0 2 0 0 16 3
708 199
708 283
575 283
1 0 4 0 0 8320 0 3 0 0 17 3
671 200
671 272
555 272
1 0 5 0 0 8320 0 4 0 0 18 3
636 200
636 266
534 266
1 0 6 0 0 8320 0 5 0 0 19 3
600 200
600 259
513 259
1 0 7 0 0 8320 0 6 0 0 9 4
293 203
293 296
401 296
401 285
1 0 8 0 0 8320 0 7 0 0 7 2
372 203
372 258
3 1 8 0 0 128 0 8 15 0 0 2
353 258
417 258
2 0 9 0 0 4096 0 15 0 0 14 2
417 276
406 276
3 1 7 0 0 128 0 15 1 0 0 2
417 285
397 285
10 0 2 0 0 4096 0 15 0 0 12 2
481 285
500 285
9 0 2 0 0 0 0 15 0 0 12 2
481 276
500 276
8 1 2 0 0 8320 0 15 13 0 0 3
481 267
500 267
500 370
7 0 9 0 0 12288 0 15 0 0 14 4
481 258
485 258
485 231
406 231
6 1 9 0 0 8320 0 15 14 0 0 3
411 330
406 330
406 226
5 0 3 0 0 128 0 15 0 0 16 5
417 312
394 312
394 345
488 345
488 330
1 14 3 0 0 0 0 9 15 0 0 3
575 248
575 330
481 330
1 13 4 0 0 128 0 10 15 0 0 3
555 248
555 321
481 321
1 12 5 0 0 128 0 11 15 0 0 3
534 248
534 312
481 312
1 11 6 0 0 128 0 12 15 0 0 3
513 248
513 303
481 303
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
