CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 200 10
216 97 1918 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
13 C:\CM\BOM.DAT
0 7
5 4 0.235825 0.500000
426 217 567 338
177209362 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 171 278 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
1 d
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
41714.8 0
0
13 Logic Switch~
5 170 232 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -17 8 -9
1 c
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
41714.8 1
0
13 Logic Switch~
5 171 177 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
1 b
-4 -27 3 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
41714.8 2
0
13 Logic Switch~
5 169 122 0 1 11
0 6
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 a
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
41714.8 3
0
2 +V
167 513 240 0 1 3
0 2
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.8956e-315 0
0
6 74LS74
17 502 158 0 12 25
0 3 5 2 2 13 14 15 16 4
5 17 18
0
0 0 5104 0
6 74LS74
-20 -70 22 -62
2 U3
-7 -61 7 -53
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 3 2 4 1 11 12 10 13 5
6 9 8 3 2 4 1 11 12 10
13 5 6 9 8 12847868
65 0 0 512 1 1 0 0
1 U
5572 0 0
2
41714.8 4
0
14 Logic Display~
6 581 141 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
41714.8 5
0
10 2-In NAND~
219 323 141 0 3 22
0 9 10 12
0
0 0 624 0
4 4011
-7 -24 21 -16
6 NAND2A
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 5 0
1 U
7361 0 0
2
5.8956e-315 5.26354e-315
0
5 4023~
219 291 234 0 4 22
0 8 7 6 11
0
0 0 624 0
4 4023
-14 -28 14 -20
5 NAND3
-19 -25 16 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 26
65 0 0 0 3 2 4 0
1 U
4747 0 0
2
5.8956e-315 5.30499e-315
0
10 2-In NAND~
219 396 194 0 3 22
0 12 11 3
0
0 0 624 0
4 4011
-7 -24 21 -16
6 NAND2B
-22 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 5 0
1 U
972 0 0
2
41714.8 6
0
9 Inverter~
13 236 132 0 2 22
0 6 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 5 1 0
1 U
3472 0 0
2
41714.8 7
0
14 Logic Display~
6 466 249 0 1 2
10 3
0
0 0 53856 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
41714.8 8
0
14
4 1 2 0 0 4224 0 6 5 0 0 6
464 149
464 227
503 227
503 262
513 262
513 249
3 4 2 0 0 0 0 6 6 0 0 2
464 140
464 149
0 1 3 0 0 4224 0 0 12 4 0 3
449 122
449 235
466 235
1 3 3 0 0 0 0 6 10 0 0 3
470 122
423 122
423 194
1 9 4 0 0 8320 0 7 6 0 0 3
565 145
565 131
534 131
2 10 5 0 0 12416 0 6 6 0 0 6
470 131
460 131
460 85
548 85
548 140
540 140
0 3 6 0 0 4224 0 0 9 11 0 3
194 122
194 243
267 243
1 2 7 0 0 8320 0 2 9 0 0 3
182 232
182 234
267 234
1 1 8 0 0 4224 0 3 9 0 0 4
183 177
259 177
259 225
267 225
2 1 9 0 0 4224 0 11 8 0 0 2
257 132
299 132
1 1 6 0 0 0 0 4 11 0 0 4
181 122
194 122
194 132
221 132
1 2 10 0 0 8320 0 1 8 0 0 4
183 278
226 278
226 150
299 150
4 2 11 0 0 4224 0 9 10 0 0 4
318 234
357 234
357 203
372 203
1 3 12 0 0 8320 0 10 8 0 0 4
372 185
357 185
357 141
350 141
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
