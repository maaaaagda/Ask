CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 429 285 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89559e-315 0
0
13 Logic Switch~
5 436 228 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89559e-315 5.26354e-315
0
13 Logic Switch~
5 439 183 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89559e-315 5.30499e-315
0
7 Ground~
168 404 316 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
5.89559e-315 5.32571e-315
0
9 Inverter~
13 539 306 0 2 22
0 9 10
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8157 0 0
2
5.89559e-315 5.34643e-315
0
7 74LS194
49 489 249 0 14 29
0 5 4 2 11 10 3 12 13 14
15 6 7 8 9
0
0 0 4848 0
6 74F194
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
5572 0 0
2
5.89559e-315 5.3568e-315
0
14 Logic Display~
6 608 215 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89559e-315 5.36716e-315
0
14 Logic Display~
6 583 215 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.89559e-315 5.37752e-315
0
14 Logic Display~
6 560 215 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89559e-315 5.38788e-315
0
14 Logic Display~
6 537 216 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89559e-315 5.39306e-315
0
10
6 1 3 0 0 4224 0 6 1 0 0 2
451 285
441 285
2 1 4 0 0 4224 0 6 2 0 0 3
457 231
448 231
448 228
3 1 2 0 0 8320 0 6 4 0 0 3
457 240
404 240
404 310
1 1 5 0 0 8320 0 6 3 0 0 3
457 213
451 213
451 183
11 1 6 0 0 8320 0 6 10 0 0 3
521 258
537 258
537 234
12 1 7 0 0 4224 0 6 9 0 0 3
521 267
560 267
560 233
13 1 8 0 0 4224 0 6 8 0 0 3
521 276
583 276
583 233
0 1 9 0 0 4224 0 0 7 9 0 3
525 285
608 285
608 233
14 1 9 0 0 0 0 6 5 0 0 4
521 285
525 285
525 306
524 306
5 2 10 0 0 12416 0 6 5 0 0 5
457 267
452 267
452 323
560 323
560 306
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
