CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 120 1 200 10
176 79 1364 538
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.268025 0.500000
176 547 1364 717
9437202 0
0
6 Title:
5 Name:
0
0
0
17
13 Logic Switch~
5 359 296 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7121 0 0
2
40240.6 0
0
5 SCOPE
12 712 169 0 1 11
0 5
0
0 0 57584 0
2 Q0
-8 -4 6 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4484 0 0
2
40240.6 0
0
5 SCOPE
12 677 169 0 1 11
0 6
0
0 0 57584 0
2 Q1
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5996 0 0
2
40240.6 0
0
5 SCOPE
12 641 169 0 1 11
0 7
0
0 0 57584 0
2 Q2
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7804 0 0
2
40240.6 0
0
5 SCOPE
12 605 169 0 1 11
0 8
0
0 0 57584 0
2 Q3
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5523 0 0
2
40240.6 0
0
5 SCOPE
12 434 394 0 1 11
0 3
0
0 0 57584 180
3 DSL
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3330 0 0
2
40240.6 0
0
5 SCOPE
12 382 394 0 1 11
0 4
0
0 0 57584 180
3 CLR
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3465 0 0
2
40240.6 0
0
5 SCOPE
12 376 166 0 1 11
0 9
0
0 0 57584 0
3 CLK
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8396 0 0
2
40240.6 0
0
14 Logic Display~
6 577 209 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
5.89467e-315 0
0
7 Pulser~
4 340 233 0 10 12
0 11 12 9 13 0 0 2 2 1
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7849 0 0
2
40240.6 1
0
7 Ground~
168 403 356 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6343 0 0
2
40240.6 2
0
14 Logic Display~
6 555 209 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
40240.6 3
0
14 Logic Display~
6 534 209 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
40240.6 4
0
14 Logic Display~
6 512 209 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
40240.6 5
0
9 Inverter~
13 454 326 0 2 22
0 5 3
0
0 0 624 512
6 74LS04
-21 -19 21 -11
3 U2A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7207 0 0
2
40240.6 6
0
2 +V
167 407 176 0 1 3
0 10
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4459 0 0
2
40240.6 7
0
7 74LS194
49 458 260 0 14 29
0 9 10 2 14 3 4 15 16 17
18 8 7 6 5
0
0 0 4848 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
3760 0 0
2
40240.6 8
0
17
1 0 3 0 0 4224 0 6 0 0 17 2
432 388
432 326
0 1 4 0 0 4224 0 0 7 8 0 2
380 296
380 388
1 0 5 0 0 8320 0 2 0 0 11 3
712 181
712 272
577 272
1 0 6 0 0 8320 0 3 0 0 14 3
677 181
677 259
555 259
1 0 7 0 0 8320 0 4 0 0 15 3
641 181
641 247
534 247
1 0 8 0 0 8320 0 5 0 0 16 3
605 181
605 235
512 235
1 0 9 0 0 4112 0 8 0 0 9 2
376 178
376 224
1 6 4 0 0 128 0 1 17 0 0 2
371 296
420 296
3 1 9 0 0 4224 0 10 17 0 0 2
364 224
426 224
0 1 5 0 0 0 0 0 15 11 0 3
496 296
496 326
475 326
14 1 5 0 0 128 0 17 9 0 0 3
490 296
577 296
577 227
3 1 2 0 0 8320 0 17 11 0 0 3
426 251
403 251
403 350
2 1 10 0 0 8320 0 17 16 0 0 3
426 242
407 242
407 185
13 1 6 0 0 128 0 17 12 0 0 3
490 287
555 287
555 227
1 12 7 0 0 128 0 13 17 0 0 3
534 227
534 278
490 278
11 1 8 0 0 128 0 17 14 0 0 3
490 269
512 269
512 227
2 5 3 0 0 128 0 15 17 0 0 4
439 326
416 326
416 278
426 278
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
