CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
230 80 30 110 10
241 79 1438 849
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
241 79 1503 849
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 489 644 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8885 0 0
2
41338.8 0
0
13 Logic Switch~
5 490 579 0 1 11
0 7
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3780 0 0
2
41338.8 0
0
13 Logic Switch~
5 497 500 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9265 0 0
2
5.89606e-315 0
0
13 Logic Switch~
5 522 320 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9442 0 0
2
5.89606e-315 0
0
13 Logic Switch~
5 667 427 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
41338.8 0
0
13 Logic Switch~
5 696 427 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9968 0 0
2
41338.8 1
0
13 Logic Switch~
5 721 427 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9281 0 0
2
41338.8 2
0
9 Inverter~
13 554 537 0 2 22
0 8 9
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
8464 0 0
2
41338.8 0
0
9 Inverter~
13 554 579 0 2 22
0 7 10
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4B
-12 -19 9 -11
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
7168 0 0
2
41338.8 0
0
9 Inverter~
13 553 500 0 2 22
0 11 12
0
0 0 624 0
5 74F04
-18 -19 17 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3171 0 0
2
41338.8 0
0
10 3-In NAND~
219 718 570 0 4 22
0 5 6 4 3
0
0 0 624 0
5 74F10
-18 -28 17 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 2 0
1 U
4139 0 0
2
41338.8 0
0
10 2-In NAND~
219 629 635 0 3 22
0 7 8 4
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6435 0 0
2
41338.8 0
0
10 2-In NAND~
219 630 570 0 3 22
0 11 10 6
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5283 0 0
2
41338.8 0
0
10 2-In NAND~
219 631 509 0 3 22
0 12 9 5
0
0 0 624 0
5 74F37
-10 -24 25 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6874 0 0
2
41338.8 0
0
14 Logic Display~
6 759 545 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
5.89606e-315 0
0
14 Logic Display~
6 756 357 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
41338.8 3
0
7 Ground~
168 588 402 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
969 0 0
2
41338.8 4
0
7 74LS151
20 639 347 0 14 29
0 13 2 13 13 13 13 2 13 2
14 15 16 17 2
0
0 0 4848 0
6 74F151
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 0 1 0 0 0
1 U
8402 0 0
2
41338.8 5
0
27
4 1 3 0 0 4224 0 11 15 0 0 3
745 570
759 570
759 563
3 3 4 0 0 8320 0 12 11 0 0 4
656 635
691 635
691 579
694 579
3 1 5 0 0 8320 0 14 11 0 0 4
658 509
691 509
691 561
694 561
3 2 6 0 0 4224 0 13 11 0 0 2
657 570
694 570
0 1 7 0 0 8320 0 0 12 10 0 3
534 579
534 626
605 626
0 2 8 0 0 4096 0 0 12 7 0 2
505 644
605 644
1 1 8 0 0 8320 0 8 1 0 0 4
539 537
505 537
505 644
501 644
2 2 9 0 0 8320 0 8 14 0 0 4
575 537
592 537
592 518
607 518
2 2 10 0 0 4224 0 9 13 0 0 2
575 579
606 579
1 1 7 0 0 0 0 2 9 0 0 2
502 579
539 579
0 1 11 0 0 8336 0 0 13 13 0 3
538 500
538 561
606 561
2 1 12 0 0 4224 0 10 14 0 0 2
574 500
607 500
1 1 11 0 0 0 0 3 10 0 0 2
509 500
538 500
4 0 13 0 0 4224 0 18 0 0 21 2
607 347
534 347
5 0 13 0 0 0 0 18 0 0 21 2
607 356
534 356
7 0 2 0 0 4096 0 18 0 0 23 2
607 374
588 374
2 0 2 0 0 0 0 18 0 0 23 2
607 329
588 329
1 1 13 0 0 128 0 18 4 0 0 2
607 320
534 320
3 0 13 0 0 0 0 18 0 0 21 2
607 338
534 338
6 0 13 0 0 0 0 18 0 0 21 2
607 365
534 365
8 1 13 0 0 0 0 18 4 0 0 3
607 383
534 383
534 320
14 1 2 0 0 8192 0 18 17 0 0 3
677 383
677 396
588 396
9 1 2 0 0 16512 0 18 17 0 0 5
677 320
683 320
683 282
588 282
588 396
10 1 14 0 0 8320 0 18 5 0 0 4
671 329
680 329
680 427
679 427
11 1 15 0 0 8320 0 18 6 0 0 3
671 338
708 338
708 427
12 1 16 0 0 8320 0 18 7 0 0 3
671 347
733 347
733 427
1 13 17 0 0 8320 0 16 18 0 0 3
756 375
756 374
671 374
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
