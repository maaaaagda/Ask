CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 170 1 240 10
176 79 1364 558
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 2 0.235110 0.500000
176 567 1364 717
42991634 0
0
6 Title:
5 Name:
0
0
0
15
5 SCOPE
12 712 209 0 1 11
0 4
0
0 0 57584 0
2 Q0
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9592 0 0
2
40240.6 0
0
5 SCOPE
12 677 209 0 1 11
0 5
0
0 0 57584 0
2 Q1
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
8748 0 0
2
40240.6 0
0
5 SCOPE
12 641 209 0 1 11
0 6
0
0 0 57584 0
2 Q2
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
7168 0 0
2
40240.6 0
0
5 SCOPE
12 606 209 0 1 11
0 7
0
0 0 57584 0
2 Q3
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
631 0 0
2
40240.6 0
0
5 SCOPE
12 351 321 0 1 11
0 3
0
0 0 57584 0
3 DSL
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
9466 0 0
2
40240.6 0
0
5 SCOPE
12 370 170 0 1 11
0 8
0
0 0 57584 0
3 CLK
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3266 0 0
2
40240.6 0
0
14 Logic Display~
6 578 242 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7693 0 0
2
5.89467e-315 0
0
14 Logic Display~
6 556 242 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3723 0 0
2
5.89467e-315 0
0
14 Logic Display~
6 534 242 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3440 0 0
2
5.89467e-315 0
0
7 Ground~
168 391 359 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6263 0 0
2
40240.6 0
0
7 Pulser~
4 335 237 0 10 12
0 10 11 8 12 0 0 2 2 2
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4900 0 0
2
40240.6 1
0
2 +V
167 403 190 0 1 3
0 9
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8783 0 0
2
40240.6 2
0
14 Logic Display~
6 513 242 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
40240.6 3
0
10 3-In NAND~
219 448 338 0 4 22
0 7 6 5 3
0
0 0 624 512
6 74LS10
-21 -28 21 -20
3 U2A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
3215 0 0
2
40240.6 4
0
7 74LS194
49 457 264 0 14 29
0 8 9 2 13 3 9 14 15 16
17 7 6 5 4
0
0 0 4848 0
7 74LS194
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 11 10 9 2 7 1 6 5 4
3 12 13 14 15 11 10 9 2 7
1 6 5 4 3 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
7903 0 0
2
40240.6 5
0
18
0 1 3 0 0 4240 0 0 5 14 0 3
415 338
351 338
351 333
1 0 4 0 0 8320 0 1 0 0 10 3
712 221
712 289
578 289
1 0 5 0 0 8320 0 2 0 0 11 3
677 221
677 280
556 280
1 0 6 0 0 8320 0 3 0 0 12 3
641 221
641 274
534 274
1 0 7 0 0 8320 0 4 0 0 13 3
606 221
606 266
513 266
1 0 8 0 0 4096 0 6 0 0 18 2
370 182
370 228
0 3 5 0 0 128 0 0 14 11 0 3
555 291
555 347
474 347
0 2 6 0 0 128 0 0 14 12 0 3
534 282
534 338
474 338
0 1 7 0 0 128 0 0 14 13 0 3
512 273
512 329
474 329
14 1 4 0 0 128 0 15 7 0 0 3
489 300
578 300
578 260
13 1 5 0 0 0 0 15 8 0 0 3
489 291
556 291
556 260
12 1 6 0 0 0 0 15 9 0 0 3
489 282
534 282
534 260
11 1 7 0 0 0 0 15 13 0 0 3
489 273
513 273
513 260
5 4 3 0 0 128 0 15 14 0 0 4
425 282
415 282
415 338
423 338
2 0 9 0 0 4096 0 15 0 0 17 2
425 246
403 246
3 1 2 0 0 8320 0 15 10 0 0 3
425 255
391 255
391 353
6 1 9 0 0 8320 0 15 12 0 0 3
419 300
403 300
403 199
3 1 8 0 0 4224 0 11 15 0 0 2
359 228
425 228
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
